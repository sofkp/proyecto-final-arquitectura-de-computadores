`timescale 1ns / 1ps

module controller(input  [6:0] op,
                  input  [2:0] funct3,
                  input        funct7b5,
                  output [1:0] ResultSrc, 
                  output MemWrite, ALUSrc, RegWrite, Jump, Branch,
                  output [1:0] ImmSrc, 
                  output [2:0] ALUControl,
                  output FP, FPlw, FPsw);
  
  wire [1:0] ALUOp; 
  
  maindec md(
    .op(op), 
    .ResultSrc(ResultSrc), 
    .MemWrite(MemWrite), 
    .Branch(Branch),
    .ALUSrc(ALUSrc), 
    .RegWrite(RegWrite), 
    .Jump(Jump), 
    .ImmSrc(ImmSrc), 
    .ALUOp(ALUOp),
    .FP(FP), .FPlw(FPlw), .FPsw(FPsw)
  ); 

  aludec  ad(
    .opb5(op[5]), 
    .funct3(funct3), 
    .funct7b5(funct7b5), 
    .ALUOp(ALUOp), 
    .ALUControl(ALUControl)
  ); 

endmodule
