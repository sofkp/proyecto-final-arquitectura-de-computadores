`timescale 1ns / 1ps
module tb_falu();
    reg clk, rst, start;
    reg [31:0] op_a, op_b;
    reg [1:0] op_code;
    reg mode_fp;
    reg round_mode;
    wire [31:0] result;
    wire valid_out;
    wire [4:0] flags;

    falu aluuu (.clk(clk),.rst(rst),.start(start),.op_a(op_a),.op_b(op_b),.op_code(op_code),.mode_fp(mode_fp),
        .round_mode(round_mode),.result(result),.valid_out(valid_out),.flags(flags));

    always #5 clk = ~clk;

    initial begin
        clk = 1; rst = 1;start = 0;round_mode = 0;mode_fp = 1; op_a = 32'h00000000; op_b = 32'h00000000; op_code = 2'b11;#10 
        rst = 0;

        // 1) 5.5 (0x40B00000) / 2 (0x40000000) = 2.75 (0x40300000)
        // NO FLAG
        start=1; op_code = 2'b11;
        op_a = 32'h40B00000; op_b = 32'h40000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 2) 2.25 (0x40100000) / 5.5 (0x40B00000) = 0.4090909 (0x3ED1745D)
        // FLAG: inexact
        start=1; op_code = 2'b11;
        op_a = 32'h40100000; op_b = 32'h40B00000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 3) 1.5 (0x3FC00000) / 1.5 (0x3FC00000) = 1.0 (0x3F800000)
        // NO FLAG
        start= 1; op_code = 2'b11;
        op_a = 32'h3FC00000; op_b = 32'h3FC00000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 4) 10.0 (0x41200000) / 4.0 (0x40800000) = 2.5 (0x40200000)
        // NO FLAG
        start= 1; op_code = 2'b11;
        op_a = 32'h41200000; op_b = 32'h40800000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 4) 0 (0x00000000) / 0 (0x00000000) → NaN (0x7FC00000)
        // FLAG: invalid
        op_a = 32'h00000000; op_b = 32'h00000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 5) Inf (0x7F800000) / Inf (0x7F800000) → NaN (0x7fc00000)
        // FLAG: invalid
        op_a = 32'h7F800000; op_b = 32'h7F800000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 6) 1.0 (0x3F800000) / 0.0 (0x00000000) = +Inf (0x7F800000)
        // FLAG: div_zero
        op_a = 32'h3F800000; op_b = 32'h00000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 7) -1.0 (0xBF800000) / 0.0 (0x00000000) = -Inf (0xFF800000)
        // FLAG: div_zero
        op_a = 32'hBF800000; op_b = 32'h00000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 8) 0 (0x00000000) / 5.0 (0x40A00000) = +0 (0x00000000)
        // NO FLAG
        op_a = 32'h00000000; op_b = 32'h40A00000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 9) -0 (0X80000000) / 2.0 (0x40000000) = -0 (0x80000000)
        // NO FLAG
        op_a = 32'h80000000; op_b = 32'h40000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 10) 1.1754943e-38 (0x00800000) / 2.0 (0x40000000) = 0x?
        // FLAG: underflow + inexact
        op_a = 32'h00800000; op_b = 32'h40000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 11) 2.3509887e-38 (0x01000000) / 1e+10 (0x501502F9) = 0x?
        // FLAG: underflow + inexact
        op_a = 32'h01000000; op_b = 32'h501502F9; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 12) 3.4028234e+38 (0x7F7FFFFF) / 0.5 (0x3F000000) = +Inf (0x7F800000)
        // FLAG: overflow + inexact
        op_a = 32'h7F7FFFFF; op_b = 32'h3F000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 13) -3.4028234e+38 (0x7F7FFFFF) / 0.5 (0x3F000000) = -Inf (0xFF800000)
        // FLAG: overflow + inexact
        op_a = 32'hFF7FFFFF; op_b = 32'h3F000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 14) 1.1754943e-38 (0x00800000) / 1e+10 (0x501502F9) = 0x0....?
        // FLAG: underflow + inexact
        op_a = 32'h00800000; op_b = 32'h501502F9; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 15) 2.3509887e-38 (0x01000000) / 1e+10 (0x501502F9) = underflow
        // FLAG: underflow + inexact
        op_a = 32'h01000000; op_b = 32'h501502F9; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // MODO FP16
        mode_fp = 0;

        // 1) 6.0 (0x4600) / 2.0 (0x4000) = 3.0 (0x4200)
        // NO FLAG
        op_a = 32'h00004600; op_b = 32'h00004000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 2) 2.25 (0x4080) / 5.5 (0x4580) ≈ 0.4091 (0x368B - 0x368C)
        // FLAG: inexact
        op_a = 32'h00004080; op_b = 32'h00004580; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 3) 1.0 (0x3C00) / 1.0 (0x3C00) = 1.0 (0x3C00)
        // NO FLAG
        op_a = 32'h00003C00; op_b = 32'h00003C00; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 4) 10.0 (0x4900) / 4.0 (0x4400) = 2.5 (0x4100)
        // NO FLAG
        op_a = 32'h00004900; op_b = 32'h00004400; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 5) 0 (0x0000) / 0 (0x0000) → NaN (0x7E00)
        // FLAG: invalid
        op_a = 32'h00000000; op_b = 32'h00000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 6) +Inf (0x7C00) / +Inf (0x7C00) → NaN (0x7E00)
        // FLAG: invalid
        op_a = 32'h00007C00; op_b = 32'h00007C00; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 7) 1.0 (0x3C00) / 0.0 (0x0000) = +Inf (0x7C00)
        // FLAG: div_zero
        op_a = 32'h00003C00; op_b = 32'h00000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 8) -1.0 (0xBC00) / 0.0 (0x0000) = -Inf (0xFC00)
        // FLAG: div_zero
        op_a = 32'h0000BC00; op_b = 32'h00000000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 9) +0 (0x0000) / 5.0 (0x4500) = +0 (0x0000)
        // NO FLAG
        op_a = 32'h00000000; op_b = 32'h00004500; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 10) -0 (0x8000) / 2.0 (0x4000) = -0 (0x8000)
        // NO FLAG
        op_a = 32'h00008000; op_b = 32'h00004000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 11) Denormal pequeño: 5.97e-8 (0x0001) / 2.0 (0x4000) ≈ 0.00000002985 (0x0000)
        // FLAG: underflow + inexact
        // PROBAR
        op_a = 32'h00000001; op_b = 32'h00004000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 12) Denormal grande: 1.2e-7 (0x0002) / 1024 (0x6400) ≈ 0.0000000001 (0x0000)
        // FLAG: underflow + inexact
        op_a = 32'h00000002; op_b = 32'h00006400; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 13) Overflow: 65504 (0x7BFF) / 0.5 (0x3800) = +Inf (0x7C00)
        // FLAG: overflow + inexact
        op_a = 32'h00007BFF; op_b = 32'h00003800; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 14) Overflow: -65504 (0xFBFF) / 0.5 (0x3800) = -Inf (0xFC00)
        // FLAG: overflow + inexact
        op_a = 32'h0000FBFF; op_b = 32'h00003800; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        // 15) Underflow extremo: 6.1e-5(0x03FF)/8192(0x7000) ≈ 0.0000000074 (0x0000)
        // FLAG: underflow + inexact
        op_a = 32'h000003FF; op_b = 32'h00007000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 16) Underflow suave: 1.2e-7(0x0002)/512(0x6000) ≈ 0.00000000023(0x0000)
        // FLAG: underflow + inexact
        op_a = 32'h00000002; op_b = 32'h00006000; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        // 18) -2.75 (0xC180) / -5.5 (0xC580) ≈ 0.5 (0x3800)
        // FLAG: inexact
        op_a = 32'h0000C180; op_b = 32'h0000C580; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        $finish;
        // 32 bits

        // add ---------------------------------
        /*
        //5555.55 + 2000.2 = 75555.75 (0x479391e0) -> 7555.7495 0x45ec1dff
        start = 1; op_code = 2'b00;
        op_a = 32'h45ad9c66; op_b = 32'h44fa0666; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // +0 + -0 = +0 (0x00000000) check
        start = 1; op_code = 2'b00;
        op_a = 32'h00000000; op_b = 32'h80000000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // +Inf + (-Inf) = NaN (0x7FC00000) check
        start = 1; op_code = 3'b000;
        op_a = 32'h7F800000; op_b = 32'hFF800000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // NaN + 5.0 = NaN (0x7FC00000) check
        start = 1; op_code = 2'b00;
        op_a = 32'h7FC00000; op_b = 32'h40A00000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // 2.2e-44 (denormal) + 1 (normal) = ~1 (0x3F800000) check
        start = 1; op_code = 2'b00;
        op_a = 32'h00000010; op_b = 32'h3F800000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
       
        //1e-45 + 3e-44 = 3.1e-44 (0x00000016)
        start = 1; op_code = 2'b00;
        op_a = 32'h00000001; op_b = 32'h00000015; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10

        
        // conmutatividad (a+b == b+a) -> -292.24353 (0xc3921f2c)+ 515.4794 (0x4400deae) = 223.23587 (0x435f3c62)
        start = 1; op_code = 2'b00;
        op_a = 32'hc3921f2c; op_b = 32'h4400deae; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        op_a = 32'h4400deae; op_b = 32'hc3921f2c; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // sub ---------------------------------
        //783.57 - 285.17 = 498.4 (0x43f93333) check
        start = 1; op_code = 2'b01;
        op_a = 32'h4443e47b; op_b = 32'h438e95c3; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
       
        // Inf - Inf = NaN (0x7FC00000)
        start = 1; op_code = 3'b001;
        op_a = 32'h7F800000; op_b = 32'h7F800000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
         
         // 0.000000000000000000000000000000000000000000011 - 0.000000000000000000000000000000000000000000006 
        // denormal- denormal = 5e-45 (0x00000004)
        start = 1; op_code = 3'b001;
        op_a = 32'h00000008; op_b = 32'h00000004; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
         
        // 7.393109e19 - -7.854292e19 = 1.5247401e+20 (0x61044008)
        start = 1; op_code = 3'b001;
        op_a = 32'h60804000; op_b = 32'he0884010; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
      
        // NaN - 1024.25 = NaN
        start = 1; op_code = 3'b001;                 
        op_a = 32'h7FC00000; op_b = 32'h44800800; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
      
      
        // 1.8894078e22 - 1024.25 = 0
        start = 1; op_code = 3'b001;                 
        op_a = 32'h64800800; op_b = 32'h44800800; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10

        // mul ---------------------------------
        
        //432.5381 (0x43d844e0) * -744.2421 (0xc43a0f7f)= -321913.063874 (0xc89d2f22) 
        start = 1; op_code = 2'b10; 
        op_a = 32'h43d844e0; op_b = 32'hc43a0f7f; #20
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // +Inf * 0 = 0 
        start = 1; op_code = 3'b010;
        op_a = 32'h7F800000; op_b = 32'h00000000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // (-Inf) * (-1) = +Inf
        start = 1; op_code = 3'b010;
        op_a = 32'hFF800000; op_b = 32'hBF800000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // 4.5e-44 (denormal) * 2 = 9e-44(0x00000040) 
        start = 1; op_code = 3'b010;
        op_a = 32'h00000020; op_b = 32'h40000000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
         // 5 * NaN = NaN
        start = 1; op_code = 3'b010;
        op_a = 32'h40a00000; op_b = 32'h7FC00000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10

        // 3.587e-42 * 3.36e-43 =  0
        start = 1; op_code = 3'b010;
        op_a = 32'h00000a00; op_b = 32'h000000f0; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10 
        
        // conmutatividad (a*b == b*a) -> 515.4794 (0x4400deae) * -723.0139 (0xc434c0e4) = 372698.771364 (0xc8b5fb58)
        start = 1; op_code = 3'b010;
        op_a = 32'h4400deae; op_b = 32'hc434c0e4; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        op_a = 32'hc434c0e4; op_b = 32'h4400deae; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // div ---------------------------------
        
        // -53.166138 (0xc254aa20) / 695.80005 (0x442df334) = -0.07641008074 (0xbd9c7ce3) check
        start = 1; op_code = 2'b11;
        op_a = 32'hc254aa20; op_b = 32'h442df334; #20
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // 1 / 0  = NaN (0x7FC00000) check
        start = 1; op_code = 2'b11; // 1 / 0
        op_a = 32'h3F800000; op_b = 32'h00000000; #20
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // 1.5845633e29 / Inf = NaN (0x7FC00000)
        start = 1; op_code = 3'b011;
        op_a = 32'h70000000; op_b = 32'h7F800000; #10
        
        // 1e-45 / 3.4028235e38 = NaN
        start = 1; op_code = 3'b011;
        op_a = 32'h00000001; op_b = 32'h7f7fffff; #10
        
        // 0.00002 (0x37a7c5ac) / 5.381e-42 (0x00000f00) = NaN (0x7e00)
        start = 1; op_code = 3'b011;
        op_a = 32'h37a7c5ac; op_b = 32'h00000f00; #10
        
        // NaN * -0.00000006007076 = NaN
        start = 1; op_code = 2'b11;                  
        op_a = 32'h7FC00000; op_b = 32'hb3810040; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10

        // -1.0178848e-28 / -1.3743895e11 = 5.925e-42 0x00001084
        start = 1; op_code = 2'b11;                  
        op_a = 32'h91010840; op_b = 32'hd2000000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10

        */

        /*
        
        //16 bits

        mode_fp = 0; 

        // add ---------------------------------
        
        // 0.5 (0x3800) + 2.25 (0x4080) ≈ 2.75 (0x00004180) check
        start = 1; op_code = 2'b00;
        op_a = 32'h00003800; op_b = 32'h00004080; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // +INf (0x7C00) + 1.0 (0x3C00) = +Inf
        start = 1; op_code = 2'b00;
        op_a = 32'h00007C00; op_b = 32'h00003C00; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        // -inf (0xFC00) + 1.0 (0x3C00) = -inf
        start = 1; op_code = 2'b00;
        op_a = 32'h0000FC00; op_b = 32'h00003C00; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        //+inf (0x7C00) + -Inf (0xFC00) = NaN (0x7E00)
        start = 1; op_code = 2'b00;
        op_a = 32'h00007C00; op_b = 32'h0000FC00; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        //NaN (0x7E00) + -2.0 (0x4000) = NaN
        start = 1; op_code = 2'b00;
        op_a = 32'h00007E00; op_b = 32'h0000c000; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        // 0.00006(0x0001) + 1.0 (0x3C00)= 1.00006 (0x3C00)
        start = 1; op_code = 2'b00;
        op_a = 32'h00000001; op_b = 32'h00003C00; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        //  0.000000834465 + -5.9604645e-8 = -7.74860355e-7 0x800d
        start = 1; op_code = 2'b00;
        op_a = 32'h0000000e; op_b = 32'h00008001; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        //sub 
        
        // 0.00000017881393 (0x0003) - 0.00000011920929(0x0002) = 0 -> 0x0001
        start = 1; op_code = 2'b01;
        op_a = 32'h00000003; op_b = 32'h00000002; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        //0.0029182434  (0x19fa) - -Inf (0xFC00) = +inf (0x7c00)
        start = 1; op_code = 2'b01;                   
        op_a = 32'h000019fa; op_b = 32'h0000FC00; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        // 466.75 (0x5f4b)  -  -466.75 (0xdf4b) = 933.5 (0x634b)
        start = 1; op_code = 2'b01;
        op_a = 32'h00005f4b; op_b = 32'h0000df4b; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // 252.375 (0x5be3)  -  155.55 (0x58dc) = 96.825 (0x560d)
        start = 1; op_code = 2'b01;
        op_a = 32'h00005be3; op_b = 32'h000058dc; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        // mul
       
        // 1.75 * 2 = 3.5 (0x00004300) CHECK
        start = 1; op_code = 2'b10;
        op_a = 32'h00003f00; op_b = 32'h00004000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        //1e-5 (0x04C4) * 1e-5 (0x04C4) ≈ 1e-10 (underflow → 0x0000)
        start = 1; op_code = 2'b10;
        op_a = 32'h000004C4; op_b = 32'h000004C4; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        //inf* 2.0 = inf
        start = 1; op_code = 2'b10;
        op_a = 32'h00007C00; op_b = 32'h00004000; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
        //0.0 (0x0000) * inf (0x7C00) = NaN (0x7E00)
        start = 1; op_code = 2'b10;
        op_a = 32'h00000000; op_b = 32'h00007C00; #20;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
       
        // 8192 (0x7000) * 8192 (0x7000) = 67108864 -> overflow inf 0x7c00
        start = 1; op_code = 2'b10;                  
        op_a = 32'h00007000; op_b = 32'h00007000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
       
        
        // div 
        
        
        //6 / 2 = 3 (0x00004200) check
        start = 1; op_code = 2'b11;
        op_a = 32'h00004600; op_b = 32'h00004000; #10
        op_a = 32'h00000000; op_b = 32'h00000000; #10
        
        //1.0 / 0.0 = +Inf (0x7C00)
        start = 1; op_code = 2'b11;
        op_a = 32'h00003C00; op_b = 32'h00000000; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;

        //0.5 (0x3800) / 5.96e-8 (0x0004) = inf overflow
        start = 1; op_code = 2'b11;
        op_a = 32'h00003800; op_b = 32'h00000004; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
        
         //0.0 (0x0000) / inf (0x7C00) = NaN (0x7E00)
        start = 1; op_code = 2'b11;
        op_a = 32'h00000000; op_b = 32'h00007C00; #10;
        op_a = 32'h00000000; op_b = 32'h00000000; #10;
*/
        $finish;
    end

endmodule
